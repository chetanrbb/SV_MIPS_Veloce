//////////////////////////////////////////////////////////////////////////////////
// <alu_control.sv> - The following file generates control signals for alu.
// 
// Source: Github
// Modified by: Daksh Dharod (daksh@pdx.edu)
// Description: It calls the alu control operation. 
// 				The function parameter will store the operation to be conducted. 
// 				The aluop parameter will decide the opeation to be done directly or to be done from the funciton block.
//
// Modifications: The typedef values for different operations are modified to make the checking easy. These changes are only done for unit testing.  
//////////////////////////////////////////////////////////////////////////////////

`ifndef _alu_control
`define _alu_control


package AluCtrlSig_pkg1;
	typedef enum logic [3:0] {
		ADD = 4'd00,
		SUB = 4'd01, 
		AND = 4'd02, 
		NOR = 4'd03, 
		OR  = 4'd04, 
		SLT = 4'd05, 
		XOR = 4'd06
	} AluOp_t;
endpackage

module alu_control(
		input logic  [5:0] funct,
		input logic  [1:0] aluop,
		output logic [3:0] aluctl);

	import AluCtrlSig_pkg1::*;
	
	AluOp_t AluCtrlSig;
	
	logic [3:0] _funct;

	always_comb 
	begin
		unique case(funct[3:0])
			ADD:  _funct <= 4'd2;		// add 
			SUB:  _funct <= 4'd6;		// sub 
			OR:   _funct <= 4'd1;		// or 
			XOR:  _funct <= 4'd13;		// xor 
			NOR:  _funct <= 4'd12;		// nor 
			SLT:  _funct <= 4'd7;		// slt 
			default: _funct <= 4'd0;
		endcase
	end 

	always_comb begin
		case(aluop)
			2'd0: aluctl <= 4'd2;		/* add */
			2'd1: aluctl <= 4'd6;		/* sub */
			2'd2: aluctl <= _funct; 
			2'd3: aluctl <= 4'd2;		/* add */
			default: aluctl <= 0;   
		endcase
	end

endmodule

`endif
