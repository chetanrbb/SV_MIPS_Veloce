

///////////////////////////////////////////////////////////////////
// cpu_tb.sv - Test bench of the cpu file
//
///////////////////////////////////////////////////////////////////

module cpu_tb();

endmodule